module dcache(clk,reset,we,re,addr,wdata,rdata);
  input   clk, we,re;
  input reset;
  input[31:0]   addr, wdata;
  output[31:0]  rdata; 
  
  reg[31:0]   RAM[383:0]; 
 
  //assign rdata = re ? RAM[addr[31:0]]:0;
 
  assign rdata = re ? RAM[addr[8:0]]:0;
 
 
	always@(posedge clk or negedge reset)
	 begin
		if (~reset)
		begin
        RAM[0  ] <= 32'h2b7e1516;
        RAM[1  ] <= 32'h28aed2a6;
        RAM[2  ] <= 32'habf71588;
        RAM[3  ] <= 32'h09cf4f3c;
        RAM[4  ] <= 32'h3243f6a8;
        RAM[5  ] <= 32'h885a308d;
        RAM[6  ] <= 32'h313198a2;
        RAM[7  ] <= 32'he0370734;
        RAM[8  ] <= 32'h00000000;
        RAM[9  ] <= 32'h00000000;
        RAM[10 ] <= 32'h00000000;
        RAM[11 ] <= 32'h00000000;
        RAM[12 ] <= 32'h00000000;
        RAM[13 ] <= 32'h00000000;
        RAM[14 ] <= 32'h00000000;
        RAM[15 ] <= 32'h00000000;
        RAM[16 ] <= 32'h00000000;
        RAM[17 ] <= 32'h00000000;
        RAM[18 ] <= 32'h00000000;
        RAM[19 ] <= 32'h00000000;
        RAM[20 ] <= 32'h00000000;
        RAM[21 ] <= 32'h00000000;
        RAM[22 ] <= 32'h00000000;
        RAM[23 ] <= 32'h00000000;
        RAM[24 ] <= 32'h00000000;
		RAM[25 ] <= 32'h00000000;
        RAM[26 ] <= 32'h00000000;
        RAM[27 ] <= 32'h00000000;
        RAM[28 ] <= 32'h00000000;
        RAM[29 ] <= 32'h00000000;
        RAM[30 ] <= 32'h00000000;
        RAM[31 ] <= 32'h00000000;
        RAM[32 ] <= 32'h00000000;
        RAM[33 ] <= 32'h00000000;
        RAM[34 ] <= 32'h00000000;
        RAM[35 ] <= 32'h00000000;
        RAM[36 ] <= 32'h00000000;
        RAM[37 ] <= 32'h00000000;
        RAM[38 ] <= 32'h00000000;
        RAM[39 ] <= 32'h00000000;
        RAM[40 ] <= 32'h00000000;
        RAM[41 ] <= 32'h00000000;
        RAM[42 ] <= 32'h00000000;
        RAM[43 ] <= 32'h00000000;
        RAM[44 ] <= 32'h00000000;
        RAM[45 ] <= 32'h00000000;
        RAM[46 ] <= 32'h00000000;
        RAM[47 ] <= 32'h00000000;
        RAM[48 ] <= 32'h00000000;
        RAM[49 ] <= 32'h00000000;
        RAM[50 ] <= 32'h00000000;
        RAM[51 ] <= 32'h00000000;
        RAM[52 ] <= 32'h00000000;
        RAM[53 ] <= 32'h00000000;
        RAM[54 ] <= 32'h00000000;
        RAM[55 ] <= 32'h00000000;
        RAM[56 ] <= 32'h00000000;
        RAM[57 ] <= 32'h00000000;
        RAM[58 ] <= 32'h00000000;
        RAM[59 ] <= 32'h00000000;
        RAM[60 ] <= 32'h00000000;
        RAM[61 ] <= 32'h00000000;
        RAM[62 ] <= 32'h00000000;
        RAM[63 ] <= 32'h00000000;
        RAM[64 ] <= 32'h00000000;
        RAM[65 ] <= 32'h00000000;
        RAM[66 ] <= 32'h00000000;
        RAM[67 ] <= 32'h00000000;
        RAM[68 ] <= 32'h00000000;
        RAM[69 ] <= 32'h00000000;
        RAM[70 ] <= 32'h00000000;
        RAM[71 ] <= 32'h00000000;
        RAM[72 ] <= 32'h00000000;
        RAM[73 ] <= 32'h00000000;
        RAM[74 ] <= 32'h00000000;
        RAM[75 ] <= 32'h00000000;
        RAM[76 ] <= 32'h00000000;
        RAM[77 ] <= 32'h00000000;
        RAM[78 ] <= 32'h00000000;
        RAM[79 ] <= 32'h00000000;
        RAM[80 ] <= 32'h00000000;
        RAM[81 ] <= 32'h00000000;
        RAM[82 ] <= 32'h00000000;
        RAM[83 ] <= 32'h00000000;
        RAM[84 ] <= 32'h00000000;
        RAM[85 ] <= 32'h00000000;
        RAM[86 ] <= 32'h00000000;
        RAM[87 ] <= 32'h00000000;
        RAM[88 ] <= 32'h00000000;
        RAM[89 ] <= 32'h00000000;
        RAM[90 ] <= 32'h00000000;
        RAM[91 ] <= 32'h00000000;
        RAM[92 ] <= 32'h00000000;
        RAM[93 ] <= 32'h00000000;
        RAM[94 ] <= 32'h00000000;
        RAM[95 ] <= 32'h00000000;
        RAM[96 ] <= 32'h00000000;
        RAM[97 ] <= 32'h00000000;
        RAM[98 ] <= 32'h00000000;
        RAM[99 ] <= 32'h00000000;
        RAM[100] <= 32'h00000000;
        RAM[101] <= 32'h00000000;
        RAM[102] <= 32'h00000000;
        RAM[103] <= 32'h00000000;
        RAM[104] <= 32'h00000000;
        RAM[105] <= 32'h00000000;
        RAM[106] <= 32'h00000000;
        RAM[107] <= 32'h00000000;
        RAM[108] <= 32'h00000000;
        RAM[109] <= 32'h00000000;
        RAM[110] <= 32'h00000000;
        RAM[111] <= 32'h00000000;
        RAM[112] <= 32'h00000000;
        RAM[113] <= 32'h00000000;
        RAM[114] <= 32'h00000000;
        RAM[115] <= 32'h00000000;
        RAM[116] <= 32'h00000000;
        RAM[117] <= 32'h00000000;
        RAM[118] <= 32'h00000000;
        RAM[119] <= 32'h00000000;
        RAM[120] <= 32'h00000000;
        RAM[121] <= 32'h00000000;
        RAM[122] <= 32'h00000000;
        RAM[123] <= 32'h00000000;
        RAM[124] <= 32'h00000000;
        RAM[125] <= 32'h00000000;
        RAM[126] <= 32'h00000000;
		RAM[127] <= 32'h00000000; 		
        RAM[128] <= 32'h00000063;
        RAM[129] <= 32'h0000007c;
        RAM[130] <= 32'h00000077;
        RAM[131] <= 32'h0000007b;
        RAM[132] <= 32'h000000f2;
        RAM[133] <= 32'h0000006b;
        RAM[134] <= 32'h0000006f;
        RAM[135] <= 32'h000000c5;
        RAM[136] <= 32'h00000030;
        RAM[137] <= 32'h00000001;
        RAM[138] <= 32'h00000067;
        RAM[139] <= 32'h0000002b;
        RAM[140] <= 32'h000000fe;
        RAM[141] <= 32'h000000d7;
        RAM[142] <= 32'h000000ab;
        RAM[143] <= 32'h00000076;
        RAM[144] <= 32'h000000ca;
        RAM[145] <= 32'h00000082;
        RAM[146] <= 32'h000000c9;
        RAM[147] <= 32'h0000007d;
        RAM[148] <= 32'h000000fa;
        RAM[149] <= 32'h00000059;
        RAM[150] <= 32'h00000047;
        RAM[151] <= 32'h000000f0;
        RAM[152] <= 32'h000000ad;
        RAM[153] <= 32'h000000d4;
        RAM[154] <= 32'h000000a2;
        RAM[155] <= 32'h000000af;
        RAM[156] <= 32'h0000009c;
        RAM[157] <= 32'h000000a4;
        RAM[158] <= 32'h00000072;
        RAM[159] <= 32'h000000c0;
        RAM[160] <= 32'h000000b7;
        RAM[161] <= 32'h000000fd;
        RAM[162] <= 32'h00000093;
        RAM[163] <= 32'h00000026;
        RAM[164] <= 32'h00000036;
        RAM[165] <= 32'h0000003f;
        RAM[166] <= 32'h000000f7;
        RAM[167] <= 32'h000000cc;
        RAM[168] <= 32'h00000034;
        RAM[169] <= 32'h000000a5;
        RAM[170] <= 32'h000000e5;
        RAM[171] <= 32'h000000f1;
        RAM[172] <= 32'h00000071;
        RAM[173] <= 32'h000000d8;
        RAM[174] <= 32'h00000031;
        RAM[175] <= 32'h00000015;
        RAM[176] <= 32'h00000004;
        RAM[177] <= 32'h000000c7;
        RAM[178] <= 32'h00000023;
        RAM[179] <= 32'h000000c3;
        RAM[180] <= 32'h00000018;
        RAM[181] <= 32'h00000096;
        RAM[182] <= 32'h00000005;
        RAM[183] <= 32'h0000009a;
        RAM[184] <= 32'h00000007;
        RAM[185] <= 32'h00000012;
        RAM[186] <= 32'h00000080;
        RAM[187] <= 32'h000000e2;
        RAM[188] <= 32'h000000eb;
        RAM[189] <= 32'h00000027;
        RAM[190] <= 32'h000000b2;
        RAM[191] <= 32'h00000075;
        RAM[192] <= 32'h00000009;
        RAM[193] <= 32'h00000083;
        RAM[194] <= 32'h0000002c;
        RAM[195] <= 32'h0000001a;
        RAM[196] <= 32'h0000001b;
        RAM[197] <= 32'h0000006e;
        RAM[198] <= 32'h0000005a;
        RAM[199] <= 32'h000000a0;
        RAM[200] <= 32'h00000052;
        RAM[201] <= 32'h0000003b;
        RAM[202] <= 32'h000000d6;
        RAM[203] <= 32'h000000b3;
        RAM[204] <= 32'h00000029;
        RAM[205] <= 32'h000000e3;
        RAM[206] <= 32'h0000002f;
        RAM[207] <= 32'h00000084;
        RAM[208] <= 32'h00000053;
        RAM[209] <= 32'h000000d1;
        RAM[210] <= 32'h00000000;
        RAM[211] <= 32'h000000ed;
        RAM[212] <= 32'h00000020;
        RAM[213] <= 32'h000000fc;
        RAM[214] <= 32'h000000b1;
        RAM[215] <= 32'h0000005b;
        RAM[216] <= 32'h0000006a;
        RAM[217] <= 32'h000000cb;
        RAM[218] <= 32'h000000be;
        RAM[219] <= 32'h00000039;
        RAM[220] <= 32'h0000004a;
        RAM[221] <= 32'h0000004c;
        RAM[222] <= 32'h00000058;
        RAM[223] <= 32'h000000cf;
        RAM[224] <= 32'h000000d0;
        RAM[225] <= 32'h000000ef;
        RAM[226] <= 32'h000000aa;
        RAM[227] <= 32'h000000fb;
        RAM[228] <= 32'h00000043;
        RAM[229] <= 32'h0000004d;
        RAM[230] <= 32'h00000033;
        RAM[231] <= 32'h00000085;
        RAM[232] <= 32'h00000045;
        RAM[233] <= 32'h000000f9;
        RAM[234] <= 32'h00000002;
        RAM[235] <= 32'h0000007f;
        RAM[236] <= 32'h00000050;
        RAM[237] <= 32'h0000003c;
        RAM[238] <= 32'h0000009f;
        RAM[239] <= 32'h000000a8;
        RAM[240] <= 32'h00000051;
        RAM[241] <= 32'h000000a3;
        RAM[242] <= 32'h00000040;
        RAM[243] <= 32'h0000008f;
        RAM[244] <= 32'h00000092;
        RAM[245] <= 32'h0000009d;
        RAM[246] <= 32'h00000038;
        RAM[247] <= 32'h000000f5;
        RAM[248] <= 32'h000000bc;
        RAM[249] <= 32'h000000b6;
        RAM[250] <= 32'h000000da;
        RAM[251] <= 32'h00000021;
        RAM[252] <= 32'h00000010;
        RAM[253] <= 32'h000000ff;
        RAM[254] <= 32'h000000f3;
        RAM[255] <= 32'h000000d2;
        RAM[256] <= 32'h000000cd;
        RAM[257] <= 32'h0000000c;
        RAM[258] <= 32'h00000013;
        RAM[259] <= 32'h000000ec;
        RAM[260] <= 32'h0000005f;
        RAM[261] <= 32'h00000097;
        RAM[262] <= 32'h00000044;
        RAM[263] <= 32'h00000017;
        RAM[264] <= 32'h000000c4;
        RAM[265] <= 32'h000000a7;
        RAM[266] <= 32'h0000007e;
        RAM[267] <= 32'h0000003d;
        RAM[268] <= 32'h00000064;
        RAM[269] <= 32'h0000005d;
        RAM[270] <= 32'h00000019;
        RAM[271] <= 32'h00000073;
        RAM[272] <= 32'h00000060;
        RAM[273] <= 32'h00000081;
        RAM[274] <= 32'h0000004f;
        RAM[275] <= 32'h000000dc;
        RAM[276] <= 32'h00000022;
        RAM[277] <= 32'h0000002a;
        RAM[278] <= 32'h00000090;
        RAM[279] <= 32'h00000088;
        RAM[280] <= 32'h00000046;
        RAM[281] <= 32'h000000ee;
        RAM[282] <= 32'h000000b8;
        RAM[283] <= 32'h00000014;
        RAM[284] <= 32'h000000de;
        RAM[285] <= 32'h0000005e;
        RAM[286] <= 32'h0000000b;
        RAM[287] <= 32'h000000db;
        RAM[288] <= 32'h000000e0;
        RAM[289] <= 32'h00000032;
        RAM[290] <= 32'h0000003a;
        RAM[291] <= 32'h0000000a;
        RAM[292] <= 32'h00000049;
        RAM[293] <= 32'h00000006;
        RAM[294] <= 32'h00000024;
        RAM[295] <= 32'h0000005c;
        RAM[296] <= 32'h000000c2;
        RAM[297] <= 32'h000000d3;
        RAM[298] <= 32'h000000ac;
        RAM[299] <= 32'h00000062;
        RAM[300] <= 32'h00000091;
        RAM[301] <= 32'h00000095;
        RAM[302] <= 32'h000000e4;
        RAM[303] <= 32'h00000079;
        RAM[304] <= 32'h000000e7;
        RAM[305] <= 32'h000000c8;
        RAM[306] <= 32'h00000037;
        RAM[307] <= 32'h0000006d;
        RAM[308] <= 32'h0000008d;
        RAM[309] <= 32'h000000d5;
        RAM[310] <= 32'h0000004e;
        RAM[311] <= 32'h000000a9;
        RAM[312] <= 32'h0000006c;
        RAM[313] <= 32'h00000056;
        RAM[314] <= 32'h000000f4;
        RAM[315] <= 32'h000000ea;
        RAM[316] <= 32'h00000065;
        RAM[317] <= 32'h0000007a;
        RAM[318] <= 32'h000000ae;
        RAM[319] <= 32'h00000008;
        RAM[320] <= 32'h000000ba;
        RAM[321] <= 32'h00000078;
        RAM[322] <= 32'h00000025;
        RAM[323] <= 32'h0000002e;
        RAM[324] <= 32'h0000001c;
        RAM[325] <= 32'h000000a6;
        RAM[326] <= 32'h000000b4;
        RAM[327] <= 32'h000000c6;
        RAM[328] <= 32'h000000e8;
        RAM[329] <= 32'h000000dd;
        RAM[330] <= 32'h00000074;
        RAM[331] <= 32'h0000001f;
        RAM[332] <= 32'h0000004b;
        RAM[333] <= 32'h000000bd;
        RAM[334] <= 32'h0000008b;
        RAM[335] <= 32'h0000008a;
        RAM[336] <= 32'h00000070;
        RAM[337] <= 32'h0000003e;
        RAM[338] <= 32'h000000b5;
        RAM[339] <= 32'h00000066;
        RAM[340] <= 32'h00000048;
        RAM[341] <= 32'h00000003;
        RAM[342] <= 32'h000000f6;
        RAM[343] <= 32'h0000000e;
        RAM[344] <= 32'h00000061;
        RAM[345] <= 32'h00000035;
        RAM[346] <= 32'h00000057;
        RAM[347] <= 32'h000000b9;
        RAM[348] <= 32'h00000086;
        RAM[349] <= 32'h000000c1;
        RAM[350] <= 32'h0000001d;
        RAM[351] <= 32'h0000009e;
        RAM[352] <= 32'h000000e1;
        RAM[353] <= 32'h000000f8;
        RAM[354] <= 32'h00000098;
        RAM[355] <= 32'h00000011;
        RAM[356] <= 32'h00000069;
        RAM[357] <= 32'h000000d9;
        RAM[358] <= 32'h0000008e;
        RAM[359] <= 32'h00000094;
        RAM[360] <= 32'h0000009b;
        RAM[361] <= 32'h0000001e;
        RAM[362] <= 32'h00000087;
        RAM[363] <= 32'h000000e9;
        RAM[364] <= 32'h000000ce;
        RAM[365] <= 32'h00000055;
        RAM[366] <= 32'h00000028;
        RAM[367] <= 32'h000000df;
        RAM[368] <= 32'h0000008c;
        RAM[369] <= 32'h000000a1;
        RAM[370] <= 32'h00000089;
        RAM[371] <= 32'h0000000d;
        RAM[372] <= 32'h000000bf;
        RAM[373] <= 32'h000000e6;
        RAM[374] <= 32'h00000042;
        RAM[375] <= 32'h00000068;
        RAM[376] <= 32'h00000041;
        RAM[377] <= 32'h00000099;
        RAM[378] <= 32'h0000002d;
        RAM[379] <= 32'h0000000f;
        RAM[380] <= 32'h000000b0;
        RAM[381] <= 32'h00000054;
        RAM[382] <= 32'h000000bb;
        RAM[383] <= 32'h00000016;
		end
		else begin
			if(we)
				//RAM[addr[31:0]]<= wdata;  
				RAM[addr[8:0]]<= wdata; 
		end
	 end

	
endmodule
